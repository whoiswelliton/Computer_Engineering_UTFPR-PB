library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity hadder is
end hadder;

architecture arq of hadder is

begin


end arq;

